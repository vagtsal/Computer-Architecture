module alu(input      [31:0] a, b, 
           input      [2:0]  alucont, 
           output reg [31:0] result,
           output            zero);

  wire [31:0] b2, sum, slt;

  assign b2 = alucont[2] ? ~b:b; 
  assign sum = a + b2 + alucont[2];
  assign slt = sum[31];

  always@(*)
    case(alucont[1:0])
      2'b00: #50 result = a & b;
      2'b01: #50 result = a | b;
      2'b10: #50 result = sum;
      2'b11: #50 result = slt;
    endcase

  assign zero = (result == 32'b0);
endmodule
