library verilog;
use verilog.vl_types.all;
entity sl2_26 is
    port(
        a               : in     vl_logic_vector(25 downto 0);
        y               : out    vl_logic_vector(27 downto 0)
    );
end sl2_26;
