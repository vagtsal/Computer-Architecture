library verilog;
use verilog.vl_types.all;
entity lpm_constant4_lpm_constant_v09 is
    port(
        result          : out    vl_logic_vector(31 downto 0)
    );
end lpm_constant4_lpm_constant_v09;
